module cubic_b_spline

pub fn cubic_b_spline() {
	println('Hello World!')
}




